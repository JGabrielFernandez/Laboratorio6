LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY LECTURA_TB IS
END ENTITY;

ARCHITECTURE TB OF LECTURA_TB IS

	constant data_width : natural := 16;
	constant addr_width : natural := 12;
	constant RAM_addr_width : natural := 20;

COMPONENT Laboratorio6 IS
	PORT(
		RESET		:	IN	STD_LOGIC;
		CLK		:	IN	STD_LOGIC;
		BOTONES	: 	IN	STD_LOGIC_VECTOR(2 DOWNTO 0);				-- Boton(2): Continuar cuando error; Boton(1): Lectura; Boton(0): Escritura;
		LLAVE		:	IN	STD_LOGIC;
		
		LED_WRITE:	OUT	STD_LOGIC;
		LED_READ	:	OUT	STD_LOGIC;
		LED_ERROR:	OUT	STD_LOGIC;
		
		WE			:	OUT	STD_LOGIC;
		CE			:	OUT	STD_LOGIC;
		OE			:	OUT	STD_LOGIC;
		LB			:	OUT	STD_LOGIC;
		UB			:	OUT	STD_LOGIC;
		DATA_BUS	:	INOUT	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0);
		DATA_BUS2:	OUT	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0);
		GND		:	OUT	STD_LOGIC;
		ADDRESS	:	OUT	STD_LOGIC_VECTOR(RAM_addr_width-1 DOWNTO 0);
		
		DISP0		:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
		DISP1		:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
		DISP2		:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
		
		RAM_STATE:	OUT	STD_LOGIC_VECTOR(5 DOWNTO 0);
		TOP_STATE:	OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
		);
END COMPONENT;

COMPONENT ROM IS
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		clock			: IN STD_LOGIC  := '1';
		q				: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END COMPONENT;

SIGNAL RESET:	STD_LOGIC:='1';
SIGNAL CLK, LLAVE:	STD_LOGIC:='0';
SIGNAL LED_WRITE,LED_READ,LED_ERROR:	STD_LOGIC;
SIGNAL BOTONES	: 	STD_LOGIC_VECTOR(2 DOWNTO 0):="111";
SIGNAL ADDRESS	:	STD_LOGIC_VECTOR(RAM_addr_width-1 DOWNTO 0);
SIGNAL RADDRESS	:	STD_LOGIC_VECTOR(addr_width-1 DOWNTO 0);
SIGNAL DATA_BUS:	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0);

BEGIN
RADDRESS<=ADDRESS(addr_width-1 DOWNTO 0);
LAB6 : Laboratorio6 port map(Reset=>RESET,Clk=>CLK,Botones=>BOTONES,LED_ERROR=>LED_ERROR,LED_READ=>LED_READ,LED_WRITE=>LED_WRITE,
								WE=>OPEN,CE=>OPEN,OE=>OPEN,LB=>OPEN,UB=>OPEN,DATA_BUS=>DATA_BUS,DATA_BUS2=>OPEN,
								ADDRESS=>ADDRESS,DISP0=>OPEN,DISP1=>OPEN,DISP2=>OPEN, RAM_STATE=>OPEN,TOP_STATE=>OPEN,LLAVE=>LLAVE, GND=>OPEN);
ROM1:	ROM PORT MAP(ADDRESS=>RADDRESS,clock=>CLK,q=>DATA_BUS);
CLK <= NOT(CLK) AFTER 10ns;
ENTRADAS: PROCESS
BEGIN
WAIT UNTIL RISING_EDGE(CLK);
RESET<='0';
WAIT UNTIL RISING_EDGE(CLK);
BOTONES<="101";
WAIT UNTIL RISING_EDGE(CLK);
BOTONES<="111";
WAIT UNTIL RISING_EDGE(LED_READ);
ASSERT(FALSE) REPORT "FIN" SEVERITY FAILURE;
END PROCESS;
END TB;
