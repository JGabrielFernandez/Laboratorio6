library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Lab6_Pack is

	constant data_width : natural := 16;
	constant addr_width : natural := 20;
	 		
	constant Inicial	 : unsigned(data_width-1 downto 0) := x"0000";
	constant Final		 : unsigned(data_width-1 downto 0) := x"FFFF";









end Lab6_Pack;